LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ENVOYEUR IS
	PORT(	CLK 			: IN STD_LOGIC;
			S_OUT 		: OUT STD_LOGIC := '0';
			PARALLEL_IN : IN STD_LOGIC_VECTOR(9 DOWNTO 0));
END ENTITY ENVOYEUR;

ARCHITECTURE BEHV OF ENVOYEUR IS
BEGIN
	PROCESS(CLK) IS
	BEGIN
		IF RISING_EDGE(CLK) THEN
			S_OUT <= PARALLEL_IN(PARALLEL_IN'LENGTH-1);
		END IF;
	END PROCESS;
END ARCHITECTURE BEHV;