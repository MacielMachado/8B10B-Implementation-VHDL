LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY clockWAIT IS
	PORT ( 	CLOCK_50 : IN 	STD_LOGIC;
				newCLOCK	: OUT STD_LOGIC;
				RESET		: IN	STD_LOGIC
			);
END ENTITY clockWAIT;

ARCHITECTURE BEHV OF clockWAIT IS
	CONSTANT delay : INTEGER := 10;
	SIGNAL COUNTER : INTEGER := 0;
BEGIN
	PROCESS(CLOCK_50)
	BEGIN
	
		IF RESET = '1' THEN
			COUNTER <= 0;
			
		ELSIF RISING_EDGE(CLOCK_50) THEN
			IF COUNTER < 10 THEN
				COUNTER <= COUNTER + 1;
			ELSE
				newCLOCK <= CLOCK_50;
			END IF; -- COUNTER = 10
		END IF; -- RISING_EDGE(CLOCK_50)
		
	END PROCESS;
END ARCHITECTURE BEHV;